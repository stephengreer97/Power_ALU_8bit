// Ones Compliment

module onesCompliment(iA,A);
input A;
output iA;

nand na1(iA,A);

endmodule